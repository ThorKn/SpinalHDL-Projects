module Ulx3s (reset,
              clk25Mhz,
              tx,
              rx);

    // Input ports
    input reset;
    input clk25Mhz;
    input rx;

    // Output ports
    output tx;

    // Clock generation
    wire boardClk;
    wire boardClkLocked;

    // Instantiate a PLL to make a 10Mhz clock
    pll pll (.clkin     (clk25Mhz),
             .clkout0   (boardClk),
             .locked    (boardClkLocked));

    // Instantiate the blinky module generated by Spinal
    UartVdf uartvdf (.io_uart_txd        (tx),
                     .io_uart_rxd        (rx),
                     .clkIsLocked        (boardClkLocked),
                     .clk                (boardClk),
                     .reset              (reset));


endmodule
