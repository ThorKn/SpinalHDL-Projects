// Generator : SpinalHDL v1.3.5    git head : f0505d24810c8661a24530409359554b7cfa271a
// Date      : 24/02/2020, 11:34:25
// Component : Button


module Button (
      input   io_button,
      output  io_led);
  assign io_led = io_button;
endmodule

