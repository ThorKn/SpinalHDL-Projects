module Ulx3s (reset_in,
              clk25Mhz,
              tx,
              rx);

    // Input ports
    input reset_in;
    input clk25Mhz;
    input rx;

    // Output ports
    output tx;

    // Clock generation
    wire boardClk;

    // Instantiate a PLL to make a 10Mhz clock
    ClkDiv clkdiv (.io_clk_out     (boardClk),
                   .clk            (clk25Mhz),
                   .reset          (reset_in));

    // Instantiate the blinky module generated by Spinal
    UartVdf uartvdf (.io_uart_txd        (tx),
                     .io_uart_rxd        (rx),
                     .clk                (boardClk),
                     .reset              (reset_in));
endmodule
